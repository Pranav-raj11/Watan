1 
0 0 0 0 0 g c 1 1 47 1 
0 0 0 1 0 g c 7 1 52 1 
0 0 0 0 0 g c 15 1 11 1 
0 0 0 0 0 g c 23 1 36 1 
3 9 3 8 4 6 2 4 1 2 3 4 2 3 4 6 0 3 1 11 0 7 2 8 1 9 4 10 2 5 5 7 0 10 0 11 1 12 
11
