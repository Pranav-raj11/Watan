1 
0 1 0 0 0 g c 1 1 47 1 
0 0 0 0 0 g c 7 1 52 1 
0 0 0 0 0 g c 15 1 11 1 
0 0 0 0 0 g c 23 1 36 1 
1 10 4 6 0 12 2 8 0 3 4 11 5 7 2 8 3 9 0 3 1 10 1 4 0 6 4 9 3 4 1 11 2 2 3 5 2 5 
5
